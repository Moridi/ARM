`include "Defines.v"
module Formarding()
endmodule